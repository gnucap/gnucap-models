** NMOSFET: Benchmarking Implementation of BSIM4.8.0
.attach ./bsim480.so

** Circuit Description **
m1 2 1 0 b n1 L=0.09u W=10.0u NF=5 rgeomod=1 geomod=0
*+SA=0.5u SB=20u geomod=0 sd=0.1u
vgs 1 0 1.2 
vds 2 0 1.2 
Vb b 0 0.0 

.include modelcard.nmos

.print dc i(vds)
.dc vds 0.0 1.2 0.02 vgs 0.2 1.2 0.2 basic

.end
