DCFL inverter circuit
* from ngspice, modified

*.subckt  inv 1 2 3
*x1  1 2 3 inv
.ngspice_hfet z1 1 3 3   aload l=1u w=10u
.ngspice_hfet z2 3 2 0   adrv l=1u w=10u
*.ends

vdd  1 0 dc 2
vin  2 0 dc 0 pwl(0,0V   .5ns,0V .505ns,1V 2ns,1V)
*x1  1 2 3 inv
rload 3 0 1meg

.model adrv nhfet level=5 rd=60 rs=60 m=2.57 lambda=0.17
+ vs=1.5e5 mu=0.385 vt0=0.3 eta=1.32 sigma0=0.04
+ vsigma=0.1 vsigmat=0.3 js1s=1e-12 js1d=1e-12
+ nmax=6e15
.model aload nhfet level=5 rd=60 rs=60 m=2.57 lambda=0.17
+ vs=1.5e5 mu=0.385 vt0=-0.3 eta=1.32 sigma0=0.04
+ vsigma=0.1 vsigmat=0.3 js1s=1e-12 js1d=1e-12
+ nmax=6e15

*>.print op v(2) v(3) i(vdd)
*>.op trace iter
*>.print op vgs(z1) vgd(z1) cg(z1) cd(z1) cgd(z1)
*>.op
*>.print op gm(z1) gds(z1) ggs(z1) ggd(z1)
*>.op
*>.print op qgs(z1) cqgs(z1) qgd(z1) cqgd(z1)
*>.op
*>.print op cs(z1) p(z1)
.op
.print tran v(2) v(3) i(vdd)
.tran 0.02n 1n 

.end
