
d1 1 0 foo bar=1
.model foo sw
.op
.end
