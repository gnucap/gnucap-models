.title mos6 inverter

.width out=150

.model nmos nmos level=6 vto=0.7
.model pmos pmos level=6 vto=-0.7

.spice_mos6 Mp1 3 2 1 1 PMOS W=8e-6 L=600e-9 
.spice_mos6 Mn1 3 2 0 0 NMOS W=8e-6 L=600e-9 

.spice_mos6 Mp2 4 2 1 1 PMOS W=8e-6 L=600e-9 
.spice_mos6 Mn2 4 2 0 0 NMOS W=8e-6 L=600e-9 
R2  4 0 10k

.spice_mos6 Mp3 5 2 1 1 PMOS W=8e-6 L=600e-9 
.spice_mos6 Mn3 5 2 0 0 NMOS W=8e-6 L=600e-9 
C3  5 0 1p

.spice_mos6 Mp4 6 2 1 1 PMOS W=8e-6 L=600e-9 
R4  6 0 2.1k

.spice_mos6 Mn5 7 2 0 0 NMOS W=8e-6 L=600e-9 
R5  7 1 2.1k

vdd 1 0 5
vin 2 0 PWL (0 0, 1n 0, 3n 5, 10n 5, 12n 0, 20n 0)

.op

.print dc v(1) v(2) v(3) v(4) v(5) v(6) v(7)
.dc vin 0 5 .25

.print tran v(1) v(2) v(3) v(4) v(5) v(6) v(7)
.tran 0.1n 5n

.end
