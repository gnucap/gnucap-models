VBIC Temp test

.MODEL N1 NPN LEVEL=4 
+ IS=1e-16 IBEI=1e-18 IBEN=5e-15 IBCI=2e-17 IBCN=5e-15 ISP=1e-15 RCX=10
+ RCI=60 RBX=10 RBI=40 RE=2 RS=20 RBP=40 VEF=10 VER=4 IKF=2e-3 ITF=8e-2
+ XTF=20 IKR=2e-4 IKP=2e-4 CJE=1e-13 CJC=2e-14 CJEP=1e-13 CJCP=4e-13 VO=2
+ GAMM=2e-11 HRCF=2 QCO=1e-12 AVC1=2 AVC2=15 TF=10e-12 TR=100e-12 TD=2e-11 RTH=300

V1 1 0 1.0
VC 1 Q1_C 0.0
VB 1 Q1_B 0.0
.ngspice_vbic Q1 Q1_C Q1_B 0 N1

.OPTIONS TEMP=150
.print dc i(vc) i(vb)
.DC V1 0.2 1.2 .1

.END
