VBIC Aplac Transient Test

.MODEL N1 NPN LEVEL=4 
+ IS=1e-16 IBEI=1e-18 IBEN=5e-15 IBCI=2e-17 IBCN=5e-15 ISP=1e-15 RCX=10
+ RCI=60 RBX=10 RBI=40 RE=2 RS=20 RBP=40 VEF=10 VER=4 IKF=2e-3 ITF=8e-2
+ XTF=20 IKR=2e-4 IKP=2e-4 CJE=1e-13 CJC=2e-14 CJEP=1e-13 CJCP=4e-13 VO=2
+ GAMM=2e-11 HRCF=2 QCO=1e-12 AVC1=2 AVC2=15 TF=10e-12 TR=100e-12 TD=2e-11 RTH=300

V1 R3_P 0 5 
V2 V2_P 0 5 Pulse(0 100m 0 10n 10n 490.1n 1u)
C1 R3_N V2_P 1n  
R4 R3_N 0 100k
.ngspice_vbic Q1 R1_N R3_N Q1_E N1
R1 R3_P R1_N 100k
R2 Q1_E 0 10k
R3 R3_P R3_N 500k

.print tran v(Q1_E)
.tran 100n 10u

.END
