VBIC DiffAmp Test

.MODEL N1 NPN LEVEL=4 
+ IS=1e-16 IBEI=1e-18 IBEN=5e-15 IBCI=2e-17 IBCN=5e-15 ISP=1e-15 RCX=10
+ RCI=60 RBX=10 RBI=40 RE=2 RS=20 RBP=40 VEF=10 VER=4 IKF=2e-3 ITF=8e-2
+ XTF=20 IKR=2e-4 IKP=2e-4 CJE=1e-13 CJC=2e-14 CJEP=1e-13 CJCP=4e-13 VO=2
+ GAMM=2e-11 HRCF=2 QCO=1e-12 AVC1=2 AVC2=15 TF=10e-12 TR=100e-12 TD=2e-11 RTH=300

.MODEL P1 PNP LEVEL=4 
+ IS=1e-16 IBEI=1e-18 IBEN=5e-15 IBCI=2e-17 IBCN=5e-15 ISP=1e-15 RCX=10
+ RCI=60 RBX=10 RBI=40 RE=2 RS=20 RBP=40 VEF=10 VER=4 IKF=2e-3 ITF=8e-2
+ XTF=20 IKR=2e-4 IKP=2e-4 CJE=1e-13 CJC=2e-14 CJEP=1e-13 CJCP=4e-13 VO=2
+ GAMM=2e-11 HRCF=2 QCO=1e-12 AVC1=2 AVC2=15 TF=10e-12 TR=100e-12 TD=2e-11 RTH=300

.ngspice_vbic Q8 Q8_B Q8_B VCC P1
.ngspice_vbic Q9 Q9_B Q9_B Q8_B P1
V1 VCC 0 3.3 
V2 V2_P R3_N  AC 1 DC 0 Sine(0 10m 10Meg 0 0)
I1 VCC I1_N 10u
.ngspice_vbic Q12 Q9_B I1_N 0 N1 M=2
.ngspice_vbic Q13 Q5_B I1_N 0 N1 M=2
.ngspice_vbic Q10 Q1_E I1_N 0 N1
.ngspice_vbic Q11 I1_N I1_N 0 N1
E1 E1_P 0 Q3_C Q4_C 1
rl e1_p 0 1e6
.ngspice_vbic Q2 Q6_C R3_N Q1_E N1
R4 R3_N 0 1K
.ngspice_vbic Q3 Q3_C Q9_B Q5_C P1
.ngspice_vbic Q1 Q5_C V2_P Q1_E N1
.ngspice_vbic Q6 Q6_C Q5_B VCC P1
R1 Q3_C 0 100k
.ngspice_vbic Q7 Q5_B Q5_B VCC P1
.ngspice_vbic Q4 Q4_C Q9_B Q6_C P1
R2 Q4_C 0 100k
R3 VCC R3_N 1K
.ngspice_vbic Q5 Q5_C Q5_B VCC P1

*>.option phase=radians
*>.print op v(nodes) iter(0)
.print ac vm(e1_p) vp(e1_p)
.print tran v(e1_p)

.OP
.AC DEC 2 100k 1G

.end
doesnt seem to work
.TRAN 1n 1u 0 10n

.END
