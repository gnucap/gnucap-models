nmos n gate, linear
.width out=90
Vgs   1  0  3.236734
.spice_mos6 M1   2  1  0  4  cmosn  l= 9.u  w= 9.u  nrd= 1.  nrs= 1. 
Vds   3  0  0.01
Rds   2  3  1.
Vbs   4  0 -1.234875
.model cmosn  nmos (level=6 tox=1e-7)
.print op v(nodes) iter(0)
.op
.print op i(v*) ps(v*)
.op
.print op id(m1) is(m1) ig(m1) ib(m1) ibs(m1) ibd(m1)
.op
.print op vgs(m1) vds(m1) vbs(m1) vth(m1) vdsat(m1)
.op
.print op gmb(m1) gm(m1) gds(m1) gbd(m1) gbs(m1)
.op
.print op cgs(m1) cgd(m1) cgb(m1) cbd(m1) cbs(m1)
.op
.print op cgsovl(m1) cgdovl(m1) cgbovl(m1) cgate(m1) region(m1)
.op
.print op cgst(m1) cgdt(m1) cgbt(m1)
.op
.print op p(m1) pd(m1) ps(m1) ids(m1) idstray(m1) iderror(m1)
.op		
.print op vdm(m1) vgm(m1) vbm(m1) vsm(m1)
.op
.print op vd(m1) vg(m1) vb(m1) vs(m1)
.op
.print dc v(1) v(2) v(3) i(vds) i(rds)
.dc vgs -10 10 1
.end
