
.ngspice_bjt q1 1 2 0 foo
.model foo d
.op
.end
